module our;
    initial begin
        $display("Hello Wofdarld");
        $finish;
    end
endmodule